`define KNN_ADDR_W 3  //address width
`define KNN_WDATA_W 16 //write data width
`ifndef DATA_W
 `define DATA_W 32      //cpu data width
`endif
